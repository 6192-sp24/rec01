// Let's say we want to compute the nth fibonacci number for a fixed n.

// Sequential vs. Combinational?

module fibonacci(Empty);  // Version 1: Hardcoded number

endmodule