interface Fibonacci;
    // A way to pass in input, and a way to get the output.
endinterface

module mkFibonacci(Fibonacci);  // Version 2: Variable fibonacci

endmodule