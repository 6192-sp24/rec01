import Fibonacci::*;

// Recompile and rerun?
// make clean fibonacci_top; ./fibonacci_top

module fibonacci_top(Empty);  // Version 2.0: Variable number, our top module uses only once.

endmodule